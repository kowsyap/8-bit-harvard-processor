module mem8(clk,address,in_data,out_data,w_en,en,p_en);
//data data_mem
//256 number of 8 bit locations,8 bit data
input clk;
input[7:0] address;
input[7:0] in_data;
input en,w_en,p_en;
output [7:0] out_data;
reg[7:0] data_mem[0:255];
integer f;

initial
begin
	$readmemb("test.data", data_mem,0,255);
end
always@(*)
begin
	if(p_en==1'b1)
	begin
	f = $fopen("data_out.o");
	$fwrite(f, "time =%d\n",$time, 
	"\tdata_mem[0] = %b\n", data_mem[0],
	"\tdata_mem[1] = %b\n", data_mem[1],
	"\tdata_mem[2] = %b\n", data_mem[2],
	"\tdata_mem[3] = %b\n", data_mem[3],
	"\tdata_mem[4] = %b\n", data_mem[4],
	"\tdata_mem[5] = %b\n", data_mem[5],
	"\tdata_mem[6] = %b\n", data_mem[6],
	"\tdata_mem[7] = %b\n", data_mem[7],
	"\tdata_mem[8] = %b\n", data_mem[8],
	"\tdata_mem[9] = %b\n", data_mem[9],
	"\tdata_mem[10] = %b\n", data_mem[10],
	"\tdata_mem[11] = %b\n", data_mem[11],
	"\tdata_mem[12] = %b\n", data_mem[12],
	"\tdata_mem[13] = %b\n", data_mem[13],
	"\tdata_mem[14] = %b\n", data_mem[14],
	"\tdata_mem[15] = %b\n", data_mem[15],
	"\tdata_mem[16] = %b\n", data_mem[16],
	"\tdata_mem[17] = %b\n", data_mem[17],
	"\tdata_mem[18] = %b\n", data_mem[18],
	"\tdata_mem[19] = %b\n", data_mem[19],
	"\tdata_mem[20] = %b\n", data_mem[20],
	"\tdata_mem[21] = %b\n", data_mem[21],
	"\tdata_mem[22] = %b\n", data_mem[22],
	"\tdata_mem[23] = %b\n", data_mem[23],
	"\tdata_mem[24] = %b\n", data_mem[24],
	"\tdata_mem[25] = %b\n", data_mem[25],
	"\tdata_mem[26] = %b\n", data_mem[26],
	"\tdata_mem[27] = %b\n", data_mem[27],
	"\tdata_mem[28] = %b\n", data_mem[28],
	"\tdata_mem[29] = %b\n", data_mem[29],
	"\tdata_mem[30] = %b\n", data_mem[30],
	"\tdata_mem[31] = %b\n", data_mem[31],
	"\tdata_mem[32] = %b\n", data_mem[32],
	"\tdata_mem[33] = %b\n", data_mem[33],
	"\tdata_mem[34] = %b\n", data_mem[34],
	"\tdata_mem[35] = %b\n", data_mem[35],
	"\tdata_mem[36] = %b\n", data_mem[36],
	"\tdata_mem[37] = %b\n", data_mem[37],
	"\tdata_mem[38] = %b\n", data_mem[38],
	"\tdata_mem[39] = %b\n", data_mem[39],
	"\tdata_mem[40] = %b\n", data_mem[40],
	"\tdata_mem[41] = %b\n", data_mem[41],
	"\tdata_mem[42] = %b\n", data_mem[42],
	"\tdata_mem[43] = %b\n", data_mem[43],
	"\tdata_mem[44] = %b\n", data_mem[44],
	"\tdata_mem[45] = %b\n", data_mem[45],
	"\tdata_mem[46] = %b\n", data_mem[46],
	"\tdata_mem[47] = %b\n", data_mem[47],
	"\tdata_mem[48] = %b\n", data_mem[48],
	"\tdata_mem[49] = %b\n", data_mem[49],
	"\tdata_mem[50] = %b\n", data_mem[50],
	"\tdata_mem[51] = %b\n", data_mem[51],
	"\tdata_mem[52] = %b\n", data_mem[52],
	"\tdata_mem[53] = %b\n", data_mem[53],
	"\tdata_mem[54] = %b\n", data_mem[54],
	"\tdata_mem[55] = %b\n", data_mem[55],
	"\tdata_mem[56] = %b\n", data_mem[56],
	"\tdata_mem[57] = %b\n", data_mem[57],
	"\tdata_mem[58] = %b\n", data_mem[58],
	"\tdata_mem[59] = %b\n", data_mem[59],
	"\tdata_mem[60] = %b\n", data_mem[60],
	"\tdata_mem[61] = %b\n", data_mem[61],
	"\tdata_mem[62] = %b\n", data_mem[62],
	"\tdata_mem[63] = %b\n", data_mem[63],
	"\tdata_mem[64] = %b\n", data_mem[64],
	"\tdata_mem[65] = %b\n", data_mem[65],
	"\tdata_mem[66] = %b\n", data_mem[66],
	"\tdata_mem[67] = %b\n", data_mem[67],
	"\tdata_mem[68] = %b\n", data_mem[68],
	"\tdata_mem[69] = %b\n", data_mem[69],
	"\tdata_mem[70] = %b\n", data_mem[70],
	"\tdata_mem[71] = %b\n", data_mem[71],
	"\tdata_mem[72] = %b\n", data_mem[72],
	"\tdata_mem[73] = %b\n", data_mem[73],
	"\tdata_mem[74] = %b\n", data_mem[74],
	"\tdata_mem[75] = %b\n", data_mem[75],
	"\tdata_mem[76] = %b\n", data_mem[76],
	"\tdata_mem[77] = %b\n", data_mem[77],
	"\tdata_mem[78] = %b\n", data_mem[78],
	"\tdata_mem[79] = %b\n", data_mem[79],
	"\tdata_mem[80] = %b\n", data_mem[80],
	"\tdata_mem[81] = %b\n", data_mem[81],
	"\tdata_mem[82] = %b\n", data_mem[82],
	"\tdata_mem[83] = %b\n", data_mem[83],
	"\tdata_mem[84] = %b\n", data_mem[84],
	"\tdata_mem[85] = %b\n", data_mem[85],
	"\tdata_mem[86] = %b\n", data_mem[86],
	"\tdata_mem[87] = %b\n", data_mem[87],
	"\tdata_mem[88] = %b\n", data_mem[88],
	"\tdata_mem[89] = %b\n", data_mem[89],
	"\tdata_mem[90] = %b\n", data_mem[90],
	"\tdata_mem[91] = %b\n", data_mem[91],
	"\tdata_mem[92] = %b\n", data_mem[92],
	"\tdata_mem[93] = %b\n", data_mem[93],
	"\tdata_mem[94] = %b\n", data_mem[94],
	"\tdata_mem[95] = %b\n", data_mem[95],
	"\tdata_mem[96] = %b\n", data_mem[96],
	"\tdata_mem[97] = %b\n", data_mem[97],
	"\tdata_mem[98] = %b\n", data_mem[98],
	"\tdata_mem[99] = %b\n", data_mem[99],
	"\tdata_mem[100] = %b\n", data_mem[100],
	"\tdata_mem[101] = %b\n", data_mem[101],
	"\tdata_mem[102] = %b\n", data_mem[102],
	"\tdata_mem[103] = %b\n", data_mem[103],
	"\tdata_mem[104] = %b\n", data_mem[104],
	"\tdata_mem[105] = %b\n", data_mem[105],
	"\tdata_mem[106] = %b\n", data_mem[106],
	"\tdata_mem[107] = %b\n", data_mem[107],
	"\tdata_mem[108] = %b\n", data_mem[108],
	"\tdata_mem[109] = %b\n", data_mem[109],
	"\tdata_mem[110] = %b\n", data_mem[110],
	"\tdata_mem[111] = %b\n", data_mem[111],
	"\tdata_mem[112] = %b\n", data_mem[112],
	"\tdata_mem[113] = %b\n", data_mem[113],
	"\tdata_mem[114] = %b\n", data_mem[114],
	"\tdata_mem[115] = %b\n", data_mem[115],
	"\tdata_mem[116] = %b\n", data_mem[116],
	"\tdata_mem[117] = %b\n", data_mem[117],
	"\tdata_mem[118] = %b\n", data_mem[118],
	"\tdata_mem[119] = %b\n", data_mem[119],
	"\tdata_mem[120] = %b\n", data_mem[120],
	"\tdata_mem[121] = %b\n", data_mem[121],
	"\tdata_mem[122] = %b\n", data_mem[122],
	"\tdata_mem[123] = %b\n", data_mem[123],
	"\tdata_mem[124] = %b\n", data_mem[124],
	"\tdata_mem[125] = %b\n", data_mem[125],
	"\tdata_mem[126] = %b\n", data_mem[126],
	"\tdata_mem[127] = %b\n", data_mem[127],
	"\tdata_mem[128] = %b\n", data_mem[128],
	"\tdata_mem[129] = %b\n", data_mem[129],
	"\tdata_mem[130] = %b\n", data_mem[130],
	"\tdata_mem[131] = %b\n", data_mem[131],
	"\tdata_mem[132] = %b\n", data_mem[132],
	"\tdata_mem[133] = %b\n", data_mem[133],
	"\tdata_mem[134] = %b\n", data_mem[134],
	"\tdata_mem[135] = %b\n", data_mem[135],
	"\tdata_mem[136] = %b\n", data_mem[136],
	"\tdata_mem[137] = %b\n", data_mem[137],
	"\tdata_mem[138] = %b\n", data_mem[138],
	"\tdata_mem[139] = %b\n", data_mem[139],
	"\tdata_mem[140] = %b\n", data_mem[140],
	"\tdata_mem[141] = %b\n", data_mem[141],
	"\tdata_mem[142] = %b\n", data_mem[142],
	"\tdata_mem[143] = %b\n", data_mem[143],
	"\tdata_mem[144] = %b\n", data_mem[144],
	"\tdata_mem[145] = %b\n", data_mem[145],
	"\tdata_mem[146] = %b\n", data_mem[146],
	"\tdata_mem[147] = %b\n", data_mem[147],
	"\tdata_mem[148] = %b\n", data_mem[148],
	"\tdata_mem[149] = %b\n", data_mem[149],
	"\tdata_mem[150] = %b\n", data_mem[150],
	"\tdata_mem[151] = %b\n", data_mem[151],
	"\tdata_mem[152] = %b\n", data_mem[152],
	"\tdata_mem[153] = %b\n", data_mem[153],
	"\tdata_mem[154] = %b\n", data_mem[154],
	"\tdata_mem[155] = %b\n", data_mem[155],
	"\tdata_mem[156] = %b\n", data_mem[156],
	"\tdata_mem[157] = %b\n", data_mem[157],
	"\tdata_mem[158] = %b\n", data_mem[158],
	"\tdata_mem[159] = %b\n", data_mem[159],
	"\tdata_mem[160] = %b\n", data_mem[160],
	"\tdata_mem[161] = %b\n", data_mem[161],
	"\tdata_mem[162] = %b\n", data_mem[162],
	"\tdata_mem[163] = %b\n", data_mem[163],
	"\tdata_mem[164] = %b\n", data_mem[164],
	"\tdata_mem[165] = %b\n", data_mem[165],
	"\tdata_mem[166] = %b\n", data_mem[166],
	"\tdata_mem[167] = %b\n", data_mem[167],
	"\tdata_mem[168] = %b\n", data_mem[168],
	"\tdata_mem[169] = %b\n", data_mem[169],
	"\tdata_mem[170] = %b\n", data_mem[170],
	"\tdata_mem[171] = %b\n", data_mem[171],
	"\tdata_mem[172] = %b\n", data_mem[172],
	"\tdata_mem[173] = %b\n", data_mem[173],
	"\tdata_mem[174] = %b\n", data_mem[174],
	"\tdata_mem[175] = %b\n", data_mem[175],
	"\tdata_mem[176] = %b\n", data_mem[176],
	"\tdata_mem[177] = %b\n", data_mem[177],
	"\tdata_mem[178] = %b\n", data_mem[178],
	"\tdata_mem[179] = %b\n", data_mem[179],
	"\tdata_mem[180] = %b\n", data_mem[180],
	"\tdata_mem[181] = %b\n", data_mem[181],
	"\tdata_mem[182] = %b\n", data_mem[182],
	"\tdata_mem[183] = %b\n", data_mem[183],
	"\tdata_mem[184] = %b\n", data_mem[184],
	"\tdata_mem[185] = %b\n", data_mem[185],
	"\tdata_mem[186] = %b\n", data_mem[186],
	"\tdata_mem[187] = %b\n", data_mem[187],
	"\tdata_mem[188] = %b\n", data_mem[188],
	"\tdata_mem[189] = %b\n", data_mem[189],
	"\tdata_mem[190] = %b\n", data_mem[190],
	"\tdata_mem[191] = %b\n", data_mem[191],
	"\tdata_mem[192] = %b\n", data_mem[192],
	"\tdata_mem[193] = %b\n", data_mem[193],
	"\tdata_mem[194] = %b\n", data_mem[194],
	"\tdata_mem[195] = %b\n", data_mem[195],
	"\tdata_mem[196] = %b\n", data_mem[196],
	"\tdata_mem[197] = %b\n", data_mem[197],
	"\tdata_mem[198] = %b\n", data_mem[198],
	"\tdata_mem[199] = %b\n", data_mem[199],
	"\tdata_mem[200] = %b\n", data_mem[200],
	"\tdata_mem[201] = %b\n", data_mem[201],
	"\tdata_mem[202] = %b\n", data_mem[202],
	"\tdata_mem[203] = %b\n", data_mem[203],
	"\tdata_mem[204] = %b\n", data_mem[204],
	"\tdata_mem[205] = %b\n", data_mem[205],
	"\tdata_mem[206] = %b\n", data_mem[206],
	"\tdata_mem[207] = %b\n", data_mem[207],
	"\tdata_mem[208] = %b\n", data_mem[208],
	"\tdata_mem[209] = %b\n", data_mem[209],
	"\tdata_mem[210] = %b\n", data_mem[210],
	"\tdata_mem[211] = %b\n", data_mem[211],
	"\tdata_mem[212] = %b\n", data_mem[212],
	"\tdata_mem[213] = %b\n", data_mem[213],
	"\tdata_mem[214] = %b\n", data_mem[214],
	"\tdata_mem[215] = %b\n", data_mem[215],
	"\tdata_mem[216] = %b\n", data_mem[216],
	"\tdata_mem[217] = %b\n", data_mem[217],
	"\tdata_mem[218] = %b\n", data_mem[218],
	"\tdata_mem[219] = %b\n", data_mem[219],
	"\tdata_mem[220] = %b\n", data_mem[220],
	"\tdata_mem[221] = %b\n", data_mem[221],
	"\tdata_mem[222] = %b\n", data_mem[222],
	"\tdata_mem[223] = %b\n", data_mem[223],
	"\tdata_mem[224] = %b\n", data_mem[224],
	"\tdata_mem[225] = %b\n", data_mem[225],
	"\tdata_mem[226] = %b\n", data_mem[226],
	"\tdata_mem[227] = %b\n", data_mem[227],
	"\tdata_mem[228] = %b\n", data_mem[228],
	"\tdata_mem[229] = %b\n", data_mem[229],
	"\tdata_mem[230] = %b\n", data_mem[230],
	"\tdata_mem[231] = %b\n", data_mem[231],
	"\tdata_mem[232] = %b\n", data_mem[232],
	"\tdata_mem[233] = %b\n", data_mem[233],
	"\tdata_mem[234] = %b\n", data_mem[234],
	"\tdata_mem[235] = %b\n", data_mem[235],
	"\tdata_mem[236] = %b\n", data_mem[236],
	"\tdata_mem[237] = %b\n", data_mem[237],
	"\tdata_mem[238] = %b\n", data_mem[238],
	"\tdata_mem[239] = %b\n", data_mem[239],
	"\tdata_mem[240] = %b\n", data_mem[240],
	"\tdata_mem[241] = %b\n", data_mem[241],
	"\tdata_mem[242] = %b\n", data_mem[242],
	"\tdata_mem[243] = %b\n", data_mem[243],
	"\tdata_mem[244] = %b\n", data_mem[244],
	"\tdata_mem[245] = %b\n", data_mem[245],
	"\tdata_mem[246] = %b\n", data_mem[246],
	"\tdata_mem[247] = %b\n", data_mem[247],
	"\tdata_mem[248] = %b\n", data_mem[248],
	"\tdata_mem[249] = %b\n", data_mem[249],
	"\tdata_mem[250] = %b\n", data_mem[250],
	"\tdata_mem[251] = %b\n", data_mem[251],
	"\tdata_mem[252] = %b\n", data_mem[252],
	"\tdata_mem[253] = %b\n", data_mem[253],
	"\tdata_mem[254] = %b\n", data_mem[254],
	"\tdata_mem[255] = %b\n", data_mem[255]);
	#130;
	$fclose(f);
	end
 end
always@(posedge clk)
begin
if(w_en==1'b1)
 data_mem[address]=in_data;
end
assign out_data= (en==1'b1)? data_mem[address]:0;

endmodule